`define DATA_WIDTH 32
`define ADDR_WIDTH 32

`define MAX_DATA_RANGE 1000
`define MAX_ADDR_RANGE 1000

class template_agent extends uvm_component;
   // UVM Factory Registration
   //
   `uvm_component_utils(template_agent)

   //--------------------------------------
   //Data Members
   //--------------------------------------
endclass
